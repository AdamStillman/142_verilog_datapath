module sign_extend(in, out);
input [3:0] in;
output [15:0] out;

assign out[3:0] = in;
assign out[15] = in[3];
assign out[14] = in[3];
assign out[13] = in[3];
assign out[12] = in[3];
assign out[11] = in[3];
assign out[10] = in[3];
assign out[9] = in[3];
assign out[8] = in[3];
assign out[7] = in[3];
assign out[6] = in[3];
assign out[5] = in[3];
assign out[4] = in[3];


endmodule
