module next_address_adder(a, b, result);

input wire [15:0] a, b;

output wire[15:0] result;

assign result = a+b;


endmodule 
